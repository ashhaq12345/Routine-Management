CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
28
13 Logic Switch~
5 95 402 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 B0
-46 -1 -32 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5698 0 0
2
41811.8 0
0
13 Logic Switch~
5 93 374 0 1 11
0 20
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B1
-44 -3 -30 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5102 0 0
2
41811.8 1
0
13 Logic Switch~
5 94 342 0 1 11
0 21
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B2
-47 0 -33 8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4688 0 0
2
41811.8 2
0
13 Logic Switch~
5 91 312 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 B3
-44 -3 -30 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3689 0 0
2
41811.8 3
0
13 Logic Switch~
5 90 280 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A0
-41 -1 -27 7
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
952 0 0
2
41811.8 4
0
13 Logic Switch~
5 91 250 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-42 -3 -28 5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6913 0 0
2
41811.8 5
0
13 Logic Switch~
5 92 217 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A2
-42 -4 -28 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7615 0 0
2
41811.8 6
0
13 Logic Switch~
5 91 187 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A3
-39 -4 -25 4
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4844 0 0
2
41811.8 7
0
4 LED~
171 972 527 0 1 2
10 9
0
0 0 864 0
4 LED1
17 0 45 8
2 D8
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7939 0 0
2
5.89666e-315 0
0
4 LED~
171 889 528 0 1 2
10 8
0
0 0 864 0
4 LED1
17 0 45 8
2 D7
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3201 0 0
2
5.89666e-315 0
0
4 LED~
171 797 526 0 1 2
10 7
0
0 0 864 0
4 LED1
17 0 45 8
2 D6
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6955 0 0
2
5.89666e-315 0
0
4 LED~
171 704 522 0 1 2
10 6
0
0 0 864 0
4 LED1
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6407 0 0
2
5.89666e-315 0
0
4 LED~
171 624 522 0 1 2
10 5
0
0 0 864 0
4 LED1
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6274 0 0
2
5.89666e-315 0
0
4 LED~
171 540 518 0 1 2
10 4
0
0 0 864 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
5808 0 0
2
5.89666e-315 0
0
4 LED~
171 463 522 0 1 2
10 3
0
0 0 864 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7413 0 0
2
5.89666e-315 0
0
4 LED~
171 381 517 0 1 2
10 3
0
0 0 864 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7307 0 0
2
41811.8 8
0
9 Inverter~
13 865 143 0 2 22
0 23 27
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3664 0 0
2
41811.8 9
0
9 Inverter~
13 672 142 0 2 22
0 24 28
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9302 0 0
2
41811.8 10
0
9 Inverter~
13 459 142 0 2 22
0 25 29
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
7636 0 0
2
41811.8 11
0
9 Inverter~
13 260 137 0 2 22
0 26 30
0
0 0 608 0
5 74F04
-18 -19 17 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5208 0 0
2
41811.8 12
0
7 Ground~
168 948 227 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3951 0 0
2
41811.8 13
0
7 Ground~
168 747 218 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
423 0 0
2
41811.8 14
0
7 Ground~
168 547 216 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3608 0 0
2
41811.8 15
0
7 Ground~
168 330 209 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3819 0 0
2
41811.8 16
0
7 74LS181
132 868 247 0 22 45
0 24 23 23 24 12 12 11 10 22
21 20 19 27 2 31 32 33 34 3
4 5 6
0
0 0 4832 0
6 74F181
-21 -69 21 -61
2 U4
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
6432 0 0
2
41811.8 17
0
7 74LS181
132 672 243 0 22 45
0 25 24 24 25 15 15 14 13 22
21 20 19 28 2 35 36 37 38 12
11 10 7
0
0 0 4832 0
6 74F181
-21 -69 21 -61
2 U3
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
6846 0 0
2
41811.8 18
0
7 74LS181
132 463 238 0 22 45
0 26 25 25 26 18 18 17 16 22
21 20 19 29 2 39 40 41 42 15
14 13 8
0
0 0 4832 0
6 74F181
-21 -69 21 -61
2 U2
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
8530 0 0
2
41811.8 19
0
7 74LS181
132 261 235 0 22 45
0 2 26 26 2 2 2 2 2 22
21 20 19 30 2 43 44 45 46 18
17 16 9
0
0 0 4832 0
6 74F181
-21 -69 21 -61
2 U1
-7 -70 7 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
5702 0 0
2
41811.8 20
0
68
0 1 3 0 0 4096 0 0 16 2 0 3
463 494
381 494
381 507
19 1 3 0 0 12416 0 25 15 0 0 5
906 274
925 274
925 489
463 489
463 512
20 1 4 0 0 12416 0 25 14 0 0 5
906 283
920 283
920 495
540 495
540 508
21 1 5 0 0 12416 0 25 13 0 0 5
906 292
915 292
915 499
624 499
624 512
22 1 6 0 0 12416 0 25 12 0 0 5
906 301
910 301
910 504
704 504
704 512
22 1 7 0 0 8320 0 26 11 0 0 3
710 297
797 297
797 516
22 1 8 0 0 8320 0 27 10 0 0 9
501 292
595 292
595 508
692 508
692 547
876 547
876 510
889 510
889 518
22 1 9 0 0 12416 0 28 9 0 0 7
299 289
401 289
401 541
959 541
959 509
972 509
972 517
8 1 2 0 0 12416 0 28 24 0 0 5
223 253
174 253
174 155
330 155
330 203
7 1 2 0 0 0 0 28 24 0 0 5
223 244
179 244
179 155
330 155
330 203
6 1 2 0 0 0 0 28 24 0 0 5
223 235
184 235
184 155
330 155
330 203
5 1 2 0 0 0 0 28 24 0 0 5
223 226
189 226
189 155
330 155
330 203
21 8 10 0 0 4224 0 26 25 0 0 4
710 288
812 288
812 265
830 265
7 20 11 0 0 4224 0 25 26 0 0 4
830 256
718 256
718 279
710 279
5 6 12 0 0 4096 0 25 25 0 0 2
830 238
830 247
19 5 12 0 0 4224 0 26 25 0 0 4
710 270
822 270
822 238
830 238
21 8 13 0 0 4224 0 27 26 0 0 4
501 283
616 283
616 261
634 261
20 7 14 0 0 4224 0 27 26 0 0 4
501 274
621 274
621 252
634 252
5 6 15 0 0 4096 0 26 26 0 0 2
634 234
634 243
19 5 15 0 0 4224 0 27 26 0 0 4
501 265
626 265
626 234
634 234
21 8 16 0 0 4224 0 28 27 0 0 4
299 280
407 280
407 256
425 256
7 20 17 0 0 4224 0 27 28 0 0 4
425 247
307 247
307 271
299 271
5 6 18 0 0 4096 0 27 27 0 0 2
425 229
425 238
19 5 18 0 0 4224 0 28 27 0 0 4
299 262
417 262
417 229
425 229
12 12 19 0 0 12288 0 26 25 0 0 6
634 297
600 297
600 332
812 332
812 301
830 301
11 11 20 0 0 4096 0 25 26 0 0 6
830 292
714 292
714 322
606 322
606 288
634 288
10 10 21 0 0 12288 0 26 25 0 0 6
634 279
610 279
610 317
817 317
817 283
830 283
9 9 22 0 0 12288 0 26 25 0 0 6
634 270
630 270
630 312
822 312
822 274
830 274
12 12 19 0 0 12416 0 27 26 0 0 6
425 292
386 292
386 327
616 327
616 297
634 297
11 11 20 0 0 4096 0 26 27 0 0 6
634 288
505 288
505 317
392 317
392 283
425 283
10 10 21 0 0 12416 0 27 26 0 0 6
425 274
396 274
396 312
621 312
621 279
634 279
9 9 22 0 0 12416 0 27 26 0 0 6
425 265
421 265
421 307
626 307
626 270
634 270
12 12 19 0 0 0 0 28 27 0 0 6
223 289
184 289
184 324
402 324
402 292
425 292
11 11 20 0 0 12416 0 28 27 0 0 6
223 280
189 280
189 319
407 319
407 283
425 283
10 10 21 0 0 0 0 28 27 0 0 6
223 271
194 271
194 309
412 309
412 274
425 274
9 9 22 0 0 0 0 28 27 0 0 6
223 262
219 262
219 304
417 304
417 265
425 265
1 12 19 0 0 0 0 1 28 0 0 4
107 402
200 402
200 289
223 289
1 11 20 0 0 0 0 2 28 0 0 4
105 374
205 374
205 280
223 280
1 10 21 0 0 0 0 3 28 0 0 4
106 342
210 342
210 271
223 271
1 9 22 0 0 0 0 4 28 0 0 4
103 312
215 312
215 262
223 262
1 3 23 0 0 12416 0 8 25 0 0 6
103 187
214 187
214 160
812 160
812 220
836 220
3 4 24 0 0 12288 0 26 25 0 0 6
640 216
610 216
610 178
817 178
817 229
836 229
1 3 24 0 0 12416 0 7 26 0 0 6
104 217
194 217
194 160
616 160
616 216
640 216
3 4 25 0 0 12416 0 27 26 0 0 6
431 211
401 211
401 173
621 173
621 225
640 225
1 3 25 0 0 0 0 6 27 0 0 6
103 250
199 250
199 160
407 160
407 211
431 211
3 4 26 0 0 12416 0 28 27 0 0 6
229 208
204 208
204 165
412 165
412 220
431 220
3 1 26 0 0 0 0 28 5 0 0 4
229 208
111 208
111 280
102 280
4 1 2 0 0 0 0 28 24 0 0 5
229 217
209 217
209 170
330 170
330 203
2 13 27 0 0 8320 0 17 25 0 0 4
886 143
914 143
914 202
900 202
2 1 23 0 0 0 0 25 17 0 0 4
836 211
826 211
826 143
850 143
2 13 28 0 0 8320 0 18 26 0 0 4
693 142
718 142
718 198
704 198
2 1 24 0 0 0 0 26 18 0 0 4
640 207
630 207
630 142
657 142
2 13 29 0 0 8320 0 19 27 0 0 4
480 142
509 142
509 193
495 193
2 1 25 0 0 0 0 27 19 0 0 4
431 202
421 202
421 142
444 142
2 13 30 0 0 8320 0 20 28 0 0 4
281 137
307 137
307 190
293 190
2 1 26 0 0 0 0 28 20 0 0 4
229 199
219 199
219 137
245 137
14 1 2 0 0 0 0 25 21 0 0 3
900 211
948 211
948 221
14 1 2 0 0 0 0 26 22 0 0 3
704 207
747 207
747 212
14 1 2 0 0 0 0 27 23 0 0 3
495 202
547 202
547 210
14 1 2 0 0 0 0 28 24 0 0 3
293 199
330 199
330 203
1 4 24 0 0 0 0 25 25 0 0 4
836 202
822 202
822 229
836 229
2 3 23 0 0 0 0 25 25 0 0 2
836 211
836 220
1 4 25 0 0 0 0 26 26 0 0 4
640 198
626 198
626 225
640 225
2 3 24 0 0 0 0 26 26 0 0 2
640 207
640 216
1 4 26 0 0 0 0 27 27 0 0 4
431 193
417 193
417 220
431 220
2 3 25 0 0 0 0 27 27 0 0 2
431 202
431 211
1 4 2 0 0 0 0 28 28 0 0 4
229 190
215 190
215 217
229 217
2 3 26 0 0 0 0 28 28 0 0 2
229 199
229 208
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
